/*-
 * Copyright (c) 2014 Robert Norton
 * All rights reserved.
 *
 * This software was developed by SRI International and the University of
 * Cambridge Computer Laboratory under DARPA/AFRL contract FA8750-10-C-0237
 * ("CTSRD"), as part of the DARPA CRASH research programme.
 *
 * @BERI_LICENSE_HEADER_START@
 *
 * Licensed to BERI Open Systems C.I.C. (BERI) under one or more contributor
 * license agreements.  See the NOTICE file distributed with this work for
 * additional information regarding copyright ownership.  BERI licenses this
 * file to you under the BERI Hardware-Software License, Version 1.0 (the
 * "License"); you may not use this file except in compliance with the
 * License.  You may obtain a copy of the License at:
 *
 *   http://www.beri-open-systems.org/legal/license-1-0.txt
 *
 * Unless required by applicable law or agreed to in writing, Work distributed
 * under the License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied.  See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * @BERI_LICENSE_HEADER_END@
 *
 ******************************************************************************
 *
 * Authors: 
 *   Robert Norton <robert.norton@cl.cam.ac.uk>
 * 
 ******************************************************************************
 *
 * Description: Format of the structure used for tracing on cheri and cheri2.
 * 
 ******************************************************************************/

typedef struct {
  Bool        valid; // 1
  Bit#(4)   version; // 4
  Bit#(5)        ex; // 5
  Bit#(10)    count; // 10
  Bit#(8)      asid; // 8
  Bit#(4)  reserved; // 4
  Bit#(32)     inst; // 32
  Bit#(64)       pc; // 64
  Bit#(64)  regVal1; // 64
  Bit#(64)  regVal2; // 64
} TraceEntry deriving (Bits, Eq, FShow); // total=256
