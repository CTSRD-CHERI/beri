/*
 * Copyright (c) 2011 Jonathan Woodruff
 * All rights reserved.
 *
 * This software was developed by SRI International and the University of
 * Cambridge Computer Laboratory under DARPA/AFRL contract FA8750-10-C-0237
 * ("CTSRD"), as part of the DARPA CRASH research programme.
 *
 * @BERI_LICENSE_HEADER_START@
 *
 * Licensed to BERI Open Systems C.I.C. (BERI) under one or more contributor
 * license agreements.  See the NOTICE file distributed with this work for
 * additional information regarding copyright ownership.  BERI licenses this
 * file to you under the BERI Hardware-Software License, Version 1.0 (the
 * "License"); you may not use this file except in compliance with the
 * License.  You may obtain a copy of the License at:
 *
 *   http://www.beri-open-systems.org/legal/license-1-0.txt
 *
 * Unless required by applicable law or agreed to in writing, Work distributed
 * under the License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied.  See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * @BERI_LICENSE_HEADER_END@
 */


/*****************************************************************************

 WARNING:

 This file has been automatically generated by tools/cheri_genfiles.py
 Do not modify it by hand.

*****************************************************************************/

`define AVN_JTAG_UART_BASE	'h3f80000
`define LOOPBACK_UART_BASE	'h3f80080
`define CHERI_NET_TX	'h3f80100
`define CHERI_NET_RX	'h3f80180
`define CHERI_COUNT	'h3f80200
`define DEBUG_JTAG_UART_BASE	'h3f80280
`define CHERI_LEDS	'h3f80300
