/*****************************************************************************

 WARNING:

 This file has been automatically generated by tools/cheri_genfiles.py
 Do not modify it by hand.

*****************************************************************************/

`define AVN_JTAG_UART_BASE	'h3f80000
`define LOOPBACK_UART_BASE	'h3f80080
`define CHERI_NET_TX	'h3f80100
`define CHERI_NET_RX	'h3f80180
`define CHERI_COUNT	'h3f80200
`define DEBUG_JTAG_UART_BASE	'h3f80280
`define CHERI_LEDS	'h3f80300
