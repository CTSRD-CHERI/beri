/*-
 * Copyright (c) 2013 Jonathan Woodruff
 * All rights reserved.
 *
 * This software was developed by SRI International and the University of
 * Cambridge Computer Laboratory under DARPA/AFRL contract FA8750-10-C-0237
 * ("CTSRD"), as part of the DARPA CRASH research programme.
 *
 * @BERI_LICENSE_HEADER_START@
 *
 * Licensed to BERI Open Systems C.I.C. (BERI) under one or more contributor
 * license agreements.  See the NOTICE file distributed with this work for
 * additional information regarding copyright ownership.  BERI licenses this
 * file to you under the BERI Hardware-Software License, Version 1.0 (the
 * "License"); you may not use this file except in compliance with the
 * License.  You may obtain a copy of the License at:
 *
 *   http://www.beri-open-systems.org/legal/license-1-0.txt
 *
 * Unless required by applicable law or agreed to in writing, Work distributed
 * under the License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied.  See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * @BERI_LICENSE_HEADER_END@
 */
 (* always_ready, always_enabled *)
interface ResetBufferIfc;
  (* prefix = "" *)
  method Action resetIn(Bool reset_n_input);
  method Bool reset_n_out;
endinterface

(* synthesize, default_reset = "no_default_reset" *)
module mkResetBuffer(ResetBufferIfc);
  Reg#(Bit#(12)) count <- mkRegU;
  Wire#(Bool) start <- mkDWire(False);
  Reg#(Bool) resetReg <- mkRegU;
  
  rule countAround;
    if (count!=0) count <= count + 1;
    else if (start) count <= 1;
    else count <= 0;
  endrule
  
  rule assignResetReg;
    // Don't stay in reset state 
    resetReg <= (count == 0);
  endrule
  
  method Action resetIn(Bool reset_n_input);
    // Check the condition again because the driving circuit may be in reset.
    if (!reset_n_input) start <= True;
  endmethod
  
  method Bool reset_n_out;
    return resetReg;
  endmethod
endmodule
