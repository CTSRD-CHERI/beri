/*
* Copyright (c) 2013 Colin Rothwell
* All rights reserved.
*
* This software was developed by Colin Rothwell as part of his final year
* undergraduate project.
*
* @BERI_LICENSE_HEADER_START@
*
* Licensed to BERI Open Systems C.I.C. (BERI) under one or more contributor
* license agreements.  See the NOTICE file distributed with this work for
* additional information regarding copyright ownership.  BERI licenses this
* file to you under the BERI Hardware-Software License, Version 1.0 (the
* "License"); you may not use this file except in compliance with the
* License.  You may obtain a copy of the License at:
*
*   http://www.beri-open-systems.org/legal/license-1-0.txt
*
* Unless required by applicable law or agreed to in writing, Work distributed
* under the License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
* CONDITIONS OF ANY KIND, either express or implied.  See the License for the
* specific language governing permissions and limitations under the License.
*
* @BERI_LICENSE_HEADER_END@
*/

import CoProFPTypes::*;
import DiadicSingleMegafunctions::*;

import MegafunctionTestBench::*;

(* synthesize *)
module mkDiadicMegafunctionTests (Empty);
    let addMegafunction <- mkVerilogAddMegafunction;
    let addTb <- mkDiadicMegafunctionTestBench(addMegafunction, 7, "Add");

    let mulMegafunction <- mkVerilogMulMegafunction;
    let mulTb <- mkDiadicMegafunctionTestBench(mulMegafunction, 5, "Multiply");

    let divMegafunction <- mkVerilogDivMegafunction;
    let divTb <- mkDiadicMegafunctionTestBench(divMegafunction, 6, "Divide");

    let subMegafunction <- mkVerilogSubMegafunction;
    let subTb <- mkDiadicMegafunctionTestBench(subMegafunction, 7, "Subtract");

    rule finish(addTb.done() &&
                mulTb.done() &&
                divTb.done() &&
                subTb.done());
        $finish();
    endrule
endmodule
